module stopwatch();

endmodule 
module test_script(

);

	
endmodule 
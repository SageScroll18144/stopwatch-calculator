module main();

	//modulo keypad
	
	//modulo cronometro
	
	//modulo calculadora
	
endmodule 
module calculator();
	
endmodule 